module encoder(
    input i0,i1,i2,i3,i4,i5,i6,i7,
    output o0,o1,o2
);
    assign o0=i1|i3|i5|i7;
    assign o1=i2|i3|i6|i7;
    assign o2=i4|i5|i6|i7;
endmodule